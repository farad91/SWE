netcdf test {    // example netCDF specification in CDL
     
     dimensions:
     x = 10, y = 5;
     
     variables:
       float   z(x,y), x(x), y(y);
     
       z:units = "meters";
     
     data:
       x = -200, -100, 0, 100, 200, 300, 400, 500, 600, 700;
       y = -120, -110, -100, -90, -80;
       z =  20,21,22,23,24,25,26,27,28,29,
            30,31,32,33,34,35,36,37,38,39,
            40,41,42,43,44,45,46,47,48,49,
            50,51,52,53,54,55,56,57,58,59,
            60,61,62,63,64,65,66,67,68,69;
     }
