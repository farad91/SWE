netcdf d_test {    // example netCDF specification in CDL
     
     dimensions:
     x = 7, y = 5;
     
     variables:
       float   z(x,y), x(x), y(y);
     
       z:units = "meters";
     
     data:
       x = -100, -70, -40, -10, 20, 50, 80;
       y = -103, -102, -101, -100, -99;
       z =  01,01,01,01,01,01,01,
	        01,01,01,01,01,01,01,
	        01,01,01,01,01,01,01,
            01,01,01,01,01,01,01,
            01,01,01,01,01,01,01;
     }
