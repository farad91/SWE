netcdf test {    // example netCDF specification in CDL
     
     dimensions:
     x = 10, y = 5;
     
     variables:
       float   z(x,y), x(x), y(y);
     
       z:units = "meters";
     
     data:
       x  = 0, 10, 20, 30, 40, 50, 60, 70, 80, 90;
       y   = -140, -118, -96, -84, -52;
     }
