netcdf d_test {    // example netCDF specification in CDL
     
     dimensions:
     x = 10, y = 5;
     
     variables:
       float   z(x,y), x(x), y(y);
     
       z:units = "meters";
     
     data:
       x = -100, -70, -40, -10, 20, 50, 80;
       y = -103, -102, -101, -100, -99;
       z =  00,01,02,03,04,05,06,07,08,09,
            10,11,12,13,14,15,16,17,18,19,
            20,21,22,23,24,25,26,27,28,29,
            30,31,32,33,34,35,36,37,38,39,
            40,41,42,43,44,45,46,47,48,49;
     }
